class eth_common;
  static mailbox gen2bfm_mb=new();
  static string testcase;
endclass

