class eth_base;
  static mailbox gen2bfm_mb=new();
  static string testcase;
  static int count=8;
endclass