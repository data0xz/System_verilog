class eth_pkt_common;

  static  mailbox gen2bfm_mb=new();

endclass